interface intf;
  
  logic clk;
  logic a;
  logic b;
  logic en_i;
  logic out;
  logic en_o;
  
endinterface
