on Xilinx run cmd is ::  xrun tb.sv -uvm
