i am soukling chacha xD?
